module PontosFlutuantes(
    input logic clock ,
    input logic reset,
    input logic [0:31] op_A_in,
    input logic [0:31] op_B_in,
    output logic [0:31] data_out,
    output logic [0:3] status_out,
    output logic [0:

);
endmodule